`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:43:52 07/08/2014 
// Design Name: 
// Module Name:    back 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module back(
    input CS3,
    input [15:0] PC,
    input [15:0] IR,
    input [7:0] ALUOUT,
    output PCupdate,
    output [15:0] PCnew,
    output Rupdate,
    output [2:0] Raddr,
    output [7:0] Rdata
    );


endmodule
