`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:30:55 07/01/2014 
// Design Name: 
// Module Name:    fourtwo 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module fourtwo(
    input clk,
    input reset,
    output t1,
    output t2,
    output t3,
    output t4
    );


endmodule
